library verilog;
use verilog.vl_types.all;
entity EP4CE10 is
    generic(
        RST_CNT_LIMIT   : integer := 100;
        UART_CLK_DIVIDER: vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0);
        SENSOR_PWR_MASK_BIT: integer := 21;
        MOTOR_PWR_MASK_BIT: integer := 22;
        CAMERA_RST1_MASK_BIT: integer := 24;
        CAMERA_RST2_MASK_BIT: integer := 25;
        CAMERA_RST3_MASK_BIT: integer := 26;
        CAMERA_RST4_MASK_BIT: integer := 27;
        CAMERA_RST5_MASK_BIT: integer := 28;
        CAMERA_PWR_PULSE_TIME: integer := 5000;
        IDLE            : integer := 1;
        WAIT_FOR_PWR    : integer := 2;
        \OPEN\          : integer := 3
    );
    port(
        clkin           : in     vl_logic;
        led             : out    vl_logic;
        rs422_de_main   : out    vl_logic;
        rs422_re_n_main : out    vl_logic;
        rs422_di_main   : out    vl_logic;
        rs422_ro_main   : in     vl_logic;
        cd4514_d        : out    vl_logic_vector(3 downto 0);
        cd4514_strobe   : out    vl_logic;
        cd4514_en_n     : out    vl_logic;
        cd4514_d_1      : out    vl_logic_vector(3 downto 0);
        cd4514_strobe_1 : out    vl_logic;
        cd4514_en_n_1   : out    vl_logic;
        cd4555_d        : out    vl_logic_vector(1 downto 0);
        cd4555_en_n     : out    vl_logic;
        cd4555_d_1      : out    vl_logic_vector(1 downto 0);
        cd4555_en_n_1   : out    vl_logic;
        pre_pwr_on      : out    vl_logic;
        pre_pwr_on_1    : out    vl_logic;
        pre_pwr_on_ack  : in     vl_logic;
        camera_rst      : out    vl_logic_vector(4 downto 0);
        camera_pwr_en   : out    vl_logic_vector(4 downto 0);
        sensor_pwr_en   : out    vl_logic;
        motor_pwr_en    : out    vl_logic;
        txd_to_stm32    : out    vl_logic;
        rxd_from_stm32  : in     vl_logic
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of RST_CNT_LIMIT : constant is 1;
    attribute mti_svvh_generic_type of UART_CLK_DIVIDER : constant is 1;
    attribute mti_svvh_generic_type of SENSOR_PWR_MASK_BIT : constant is 1;
    attribute mti_svvh_generic_type of MOTOR_PWR_MASK_BIT : constant is 1;
    attribute mti_svvh_generic_type of CAMERA_RST1_MASK_BIT : constant is 1;
    attribute mti_svvh_generic_type of CAMERA_RST2_MASK_BIT : constant is 1;
    attribute mti_svvh_generic_type of CAMERA_RST3_MASK_BIT : constant is 1;
    attribute mti_svvh_generic_type of CAMERA_RST4_MASK_BIT : constant is 1;
    attribute mti_svvh_generic_type of CAMERA_RST5_MASK_BIT : constant is 1;
    attribute mti_svvh_generic_type of CAMERA_PWR_PULSE_TIME : constant is 1;
    attribute mti_svvh_generic_type of IDLE : constant is 1;
    attribute mti_svvh_generic_type of WAIT_FOR_PWR : constant is 1;
    attribute mti_svvh_generic_type of \OPEN\ : constant is 1;
end EP4CE10;
