library verilog;
use verilog.vl_types.all;
entity command_rw_main is
    generic(
        FRAME_HEAD1     : vl_logic_vector(0 to 7) := (Hi1, Hi0, Hi1, Hi0, Hi1, Hi0, Hi1, Hi0);
        FRAME_HEAD2     : vl_logic_vector(0 to 7) := (Hi0, Hi1, Hi0, Hi1, Hi0, Hi1, Hi0, Hi1);
        FRAME_HEAD3     : vl_logic_vector(0 to 7) := (Hi1, Hi1, Hi1, Hi0, Hi1, Hi0, Hi1, Hi1);
        FRAME_HEAD4     : vl_logic_vector(0 to 7) := (Hi1, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0);
        FRAME_HEAD5     : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi1, Hi1, Hi1, Hi0, Hi1);
        FRAME_HEAD6     : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi1, Hi1, Hi0, Hi1, Hi1);
        FRAME_END       : vl_logic_vector(0 to 7) := (Hi1, Hi1, Hi1, Hi0, Hi1, Hi1, Hi1, Hi1);
        IDLE            : vl_logic_vector(0 to 4) := (Hi0, Hi0, Hi0, Hi0, Hi0);
        HEAD1           : vl_logic_vector(0 to 4) := (Hi0, Hi0, Hi0, Hi0, Hi1);
        HEAD2           : vl_logic_vector(0 to 4) := (Hi0, Hi0, Hi0, Hi1, Hi0);
        HEAD3           : vl_logic_vector(0 to 4) := (Hi0, Hi0, Hi0, Hi1, Hi1);
        HEAD4           : vl_logic_vector(0 to 4) := (Hi0, Hi0, Hi1, Hi0, Hi0);
        HEAD5           : vl_logic_vector(0 to 4) := (Hi0, Hi0, Hi1, Hi0, Hi1);
        HEAD6           : vl_logic_vector(0 to 4) := (Hi0, Hi0, Hi1, Hi1, Hi0);
        COMMAND_H       : vl_logic_vector(0 to 4) := (Hi0, Hi0, Hi1, Hi1, Hi1);
        COMMAND_L       : vl_logic_vector(0 to 4) := (Hi0, Hi1, Hi0, Hi0, Hi0);
        BYTE1           : vl_logic_vector(0 to 4) := (Hi0, Hi1, Hi0, Hi0, Hi1);
        BYTE2           : vl_logic_vector(0 to 4) := (Hi0, Hi1, Hi0, Hi1, Hi0);
        BYTE3           : vl_logic_vector(0 to 4) := (Hi0, Hi1, Hi0, Hi1, Hi1);
        BYTE4           : vl_logic_vector(0 to 4) := (Hi0, Hi1, Hi1, Hi0, Hi0);
        BYTE5           : vl_logic_vector(0 to 4) := (Hi0, Hi1, Hi1, Hi0, Hi1);
        BYTE6           : vl_logic_vector(0 to 4) := (Hi0, Hi1, Hi1, Hi1, Hi0);
        CRC_H           : vl_logic_vector(0 to 4) := (Hi0, Hi1, Hi1, Hi1, Hi1);
        CRC_L           : vl_logic_vector(0 to 4) := (Hi1, Hi0, Hi0, Hi0, Hi0);
        RX_TIME_OUT_PROTECTION: integer := 100000;
        TX_GUARDING_TIME: integer := 500
    );
    port(
        uart_chip_de    : out    vl_logic;
        uart_chip_re_n  : out    vl_logic;
        uart_chip_di    : out    vl_logic;
        uart_chip_ro    : in     vl_logic;
        command_rx_ready: out    vl_logic;
        command_rx      : out    vl_logic_vector(15 downto 0);
        data_field_rx   : out    vl_logic_vector(47 downto 0);
        command_tx_over : out    vl_logic;
        command_tx_status: out    vl_logic;
        command_tx_ready: in     vl_logic;
        command_tx      : in     vl_logic_vector(15 downto 0);
        data_field_tx   : in     vl_logic_vector(47 downto 0);
        uart_clk        : in     vl_logic;
        version         : in     vl_logic_vector(31 downto 0);
        clk             : in     vl_logic;
        rst_n           : in     vl_logic
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of FRAME_HEAD1 : constant is 1;
    attribute mti_svvh_generic_type of FRAME_HEAD2 : constant is 1;
    attribute mti_svvh_generic_type of FRAME_HEAD3 : constant is 1;
    attribute mti_svvh_generic_type of FRAME_HEAD4 : constant is 1;
    attribute mti_svvh_generic_type of FRAME_HEAD5 : constant is 1;
    attribute mti_svvh_generic_type of FRAME_HEAD6 : constant is 1;
    attribute mti_svvh_generic_type of FRAME_END : constant is 1;
    attribute mti_svvh_generic_type of IDLE : constant is 1;
    attribute mti_svvh_generic_type of HEAD1 : constant is 1;
    attribute mti_svvh_generic_type of HEAD2 : constant is 1;
    attribute mti_svvh_generic_type of HEAD3 : constant is 1;
    attribute mti_svvh_generic_type of HEAD4 : constant is 1;
    attribute mti_svvh_generic_type of HEAD5 : constant is 1;
    attribute mti_svvh_generic_type of HEAD6 : constant is 1;
    attribute mti_svvh_generic_type of COMMAND_H : constant is 1;
    attribute mti_svvh_generic_type of COMMAND_L : constant is 1;
    attribute mti_svvh_generic_type of BYTE1 : constant is 1;
    attribute mti_svvh_generic_type of BYTE2 : constant is 1;
    attribute mti_svvh_generic_type of BYTE3 : constant is 1;
    attribute mti_svvh_generic_type of BYTE4 : constant is 1;
    attribute mti_svvh_generic_type of BYTE5 : constant is 1;
    attribute mti_svvh_generic_type of BYTE6 : constant is 1;
    attribute mti_svvh_generic_type of CRC_H : constant is 1;
    attribute mti_svvh_generic_type of CRC_L : constant is 1;
    attribute mti_svvh_generic_type of RX_TIME_OUT_PROTECTION : constant is 1;
    attribute mti_svvh_generic_type of TX_GUARDING_TIME : constant is 1;
end command_rw_main;
