library verilog;
use verilog.vl_types.all;
entity explosive_ctrl is
    generic(
        PRE_POWER_GUARDING_TIME: integer := 500;
        PRE_POWER_FAIL_TIME: vl_notype;
        EXPLOSION_GUARDING_TIME: vl_logic_vector(0 to 32) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi1, Hi0, Hi0, Hi1, Hi0);
        COMMAND_TYPE_EXPLODE: vl_logic_vector(0 to 15) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi1);
        COMMAND_TYPE_CANCEL: vl_logic_vector(0 to 15) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi1, Hi0);
        COMMAND_TYPE_PRE_POWER: vl_logic_vector(0 to 15) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi1, Hi1);
        IDLE            : integer := 1;
        PRE_POWER       : integer := 2;
        EXPLOSION       : integer := 3;
        OVER            : integer := 4;
        EXPLOSIVE_TIME  : integer := 1000;
        FIRE_CHANNEL1_MASK_BIT: integer := 0;
        FIRE_CHANNEL2_MASK_BIT: integer := 1;
        FIRE_CHANNEL3_MASK_BIT: integer := 2;
        FIRE_CHANNEL4_MASK_BIT: integer := 3;
        FIRE_CHANNEL5_MASK_BIT: integer := 4;
        FIRE_CHANNEL6_MASK_BIT: integer := 5;
        FIRE_CHANNEL7_MASK_BIT: integer := 6;
        FIRE_CHANNEL8_MASK_BIT: integer := 7;
        FIRE_CHANNEL9_MASK_BIT: integer := 8;
        FIRE_CHANNEL10_MASK_BIT: integer := 9;
        FIRE_CHANNEL11_MASK_BIT: integer := 10;
        FIRE_CHANNEL12_MASK_BIT: integer := 11;
        FIRE_CHANNEL13_MASK_BIT: integer := 12;
        FIRE_CHANNEL14_MASK_BIT: integer := 13;
        FIRE_CHANNEL15_MASK_BIT: integer := 14;
        FIRE_CHANNEL16_MASK_BIT: integer := 15;
        FIRE_CHANNEL17_MASK_BIT: integer := 16;
        FIRE_CHANNEL18_MASK_BIT: integer := 17;
        FIRE_CHANNEL19_MASK_BIT: integer := 18;
        FIRE_CHANNEL20_MASK_BIT: integer := 19;
        PRE_POWER_MASK_BIT: integer := 20;
        ENABLE          : vl_logic := Hi1;
        DISABLE         : vl_logic := Hi0
    );
    port(
        cd4514_d        : out    vl_logic_vector(3 downto 0);
        cd4514_strobe   : out    vl_logic;
        cd4514_en_n     : out    vl_logic;
        cd4514_d_1      : out    vl_logic_vector(3 downto 0);
        cd4514_strobe_1 : out    vl_logic;
        cd4514_en_n_1   : out    vl_logic;
        cd4555_d        : out    vl_logic_vector(1 downto 0);
        cd4555_en_n     : out    vl_logic;
        cd4555_d_1      : out    vl_logic_vector(1 downto 0);
        cd4555_en_n_1   : out    vl_logic;
        pre_pwr_on      : out    vl_logic;
        pre_pwr_on_1    : out    vl_logic;
        pre_pwr_on_ack  : in     vl_logic;
        command_ready   : in     vl_logic;
        command_type    : in     vl_logic_vector(15 downto 0);
        command_parameter: in     vl_logic_vector(31 downto 0);
        explosive_status: out    vl_logic_vector(47 downto 0);
        err_reg         : out    vl_logic_vector(7 downto 0);
        clk             : in     vl_logic;
        rst_n           : in     vl_logic
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of PRE_POWER_GUARDING_TIME : constant is 1;
    attribute mti_svvh_generic_type of PRE_POWER_FAIL_TIME : constant is 3;
    attribute mti_svvh_generic_type of EXPLOSION_GUARDING_TIME : constant is 1;
    attribute mti_svvh_generic_type of COMMAND_TYPE_EXPLODE : constant is 1;
    attribute mti_svvh_generic_type of COMMAND_TYPE_CANCEL : constant is 1;
    attribute mti_svvh_generic_type of COMMAND_TYPE_PRE_POWER : constant is 1;
    attribute mti_svvh_generic_type of IDLE : constant is 1;
    attribute mti_svvh_generic_type of PRE_POWER : constant is 1;
    attribute mti_svvh_generic_type of EXPLOSION : constant is 1;
    attribute mti_svvh_generic_type of OVER : constant is 1;
    attribute mti_svvh_generic_type of EXPLOSIVE_TIME : constant is 1;
    attribute mti_svvh_generic_type of FIRE_CHANNEL1_MASK_BIT : constant is 1;
    attribute mti_svvh_generic_type of FIRE_CHANNEL2_MASK_BIT : constant is 1;
    attribute mti_svvh_generic_type of FIRE_CHANNEL3_MASK_BIT : constant is 1;
    attribute mti_svvh_generic_type of FIRE_CHANNEL4_MASK_BIT : constant is 1;
    attribute mti_svvh_generic_type of FIRE_CHANNEL5_MASK_BIT : constant is 1;
    attribute mti_svvh_generic_type of FIRE_CHANNEL6_MASK_BIT : constant is 1;
    attribute mti_svvh_generic_type of FIRE_CHANNEL7_MASK_BIT : constant is 1;
    attribute mti_svvh_generic_type of FIRE_CHANNEL8_MASK_BIT : constant is 1;
    attribute mti_svvh_generic_type of FIRE_CHANNEL9_MASK_BIT : constant is 1;
    attribute mti_svvh_generic_type of FIRE_CHANNEL10_MASK_BIT : constant is 1;
    attribute mti_svvh_generic_type of FIRE_CHANNEL11_MASK_BIT : constant is 1;
    attribute mti_svvh_generic_type of FIRE_CHANNEL12_MASK_BIT : constant is 1;
    attribute mti_svvh_generic_type of FIRE_CHANNEL13_MASK_BIT : constant is 1;
    attribute mti_svvh_generic_type of FIRE_CHANNEL14_MASK_BIT : constant is 1;
    attribute mti_svvh_generic_type of FIRE_CHANNEL15_MASK_BIT : constant is 1;
    attribute mti_svvh_generic_type of FIRE_CHANNEL16_MASK_BIT : constant is 1;
    attribute mti_svvh_generic_type of FIRE_CHANNEL17_MASK_BIT : constant is 1;
    attribute mti_svvh_generic_type of FIRE_CHANNEL18_MASK_BIT : constant is 1;
    attribute mti_svvh_generic_type of FIRE_CHANNEL19_MASK_BIT : constant is 1;
    attribute mti_svvh_generic_type of FIRE_CHANNEL20_MASK_BIT : constant is 1;
    attribute mti_svvh_generic_type of PRE_POWER_MASK_BIT : constant is 1;
    attribute mti_svvh_generic_type of ENABLE : constant is 1;
    attribute mti_svvh_generic_type of DISABLE : constant is 1;
end explosive_ctrl;
